`timescale 1ns/1ps

module k_wctl_t1();
endmodule
